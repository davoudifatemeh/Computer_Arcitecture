<?php

$name = readline();
echo "Hello " . "$name" . "! How are you?";

php?>